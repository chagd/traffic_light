module main();

endmodule //main
